//Build a circuit with no inputs and no output that outputs a constant 1
module top_module( output one );

// Insert your code here
    assign one = 1;

endmodule
