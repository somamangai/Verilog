//Create a module that implements a NOT gate.
module top_module( input in, output out );

    assign out = !in;
endmodule
